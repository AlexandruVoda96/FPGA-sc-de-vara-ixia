module transcodor (input [6:0] points,
						 output reg [13:0] q);
	
			always@(points)
				case(points)
					  0: q=14'b10000001000000; //0
					  1: q=14'b10000001111001; //1
					  2: q=14'b10000000100100; //2
					  3: q=14'b10000000110000; //3
					  4: q=14'b10000000011001; //4
					  5: q=14'b10000000010010; //5
					  6: q=14'b10000000000010; //6
					  7: q=14'b10000001111000; //7
					  8: q=14'b10000000000000; //8
					  9: q=14'b10000000010000; //9
					  10: q=14'b11110011000000; //10
					  11: q=14'b11110011111001; //11
					  12: q=14'b11110010100100; //12
					  13: q=14'b11110010110000; //13
					  14: q=14'b11110010011001; //14
					  15: q=14'b11110010010010; //15
					  16: q=14'b11110010000010; //16
					  17: q=14'b11110011111000; //17
					  18: q=14'b11110010000000; //18
					  19: q=14'b11110010010000; //19
					  20: q=14'b01001001000000; //20
					  21: q=14'b01001001111001; //21
					  22: q=14'b01001000100100; //22
					  23: q=14'b01001000110000; //23
					  24: q=14'b01001000011001; //24
					  25: q=14'b01001000010010; //25
					  26: q=14'b01001000000010; //26
					  27: q=14'b01001001111000; //27
					  28: q=14'b01001000000000; //28
					  29: q=14'b01001000010000; //29
					  30: q=14'b01100001000000; //30
					 // 31: q=14'b01100001111001; //31
					  default:    q=14'b01100001000000;
					  
				endcase
			
endmodule