module transcodor (input [7:0] in, 
output reg[6:0] out);

always @*
case (in)
8'b01000101: out=7'b0000001; //0
8'b00010110: out=7'b1001111; //1
8'b00011110: out=7'b0010010; //2
8'b00100110: out=7'b0000110; //3
8'b00100101: out=7'b1001100; //4
8'b00101110: out=7'b0100100; //5
8'b00110110: out=7'b0100000; //6
8'b00111101: out=7'b0001111; //7
8'b00111110: out=7'b0000000; //8
8'b01000110: out=7'b0000100; //9
8'b00011100: out=7'b0001000; //a
8'b00110010: out=7'b1100000; //b
8'b00100001: out=7'b0110001; //c
8'b00100011: out=7'b1000010; //d
8'b00100100: out=7'b0110000; //e
8'b00101011: out=7'b0111000; //f
endcase
endmodule